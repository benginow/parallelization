 `timescale 1ps/1ps

 module div(input [15:0]first, input [15:0]second, output [15:0]out
    output[15:0] modulo);
    
    

 endmodule